library verilog;
use verilog.vl_types.all;
entity ee357_alu_tb is
end ee357_alu_tb;
